module RegFile(
  input         clock,
  input         reset,
  input  [4:0]  io_b_rport_0_addr,
  output [31:0] io_b_rport_0_data,
  input  [4:0]  io_b_rport_1_addr,
  output [31:0] io_b_rport_1_data,
  input         io_b_wport_0_en,
  input  [4:0]  io_b_wport_0_addr,
  input  [31:0] io_b_wport_0_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] reg_regfile_0; // @[registerFile.scala 25:26]
  reg [31:0] reg_regfile_1; // @[registerFile.scala 25:26]
  reg [31:0] reg_regfile_2; // @[registerFile.scala 25:26]
  reg [31:0] reg_regfile_3; // @[registerFile.scala 25:26]
  reg [31:0] reg_regfile_4; // @[registerFile.scala 25:26]
  reg [31:0] reg_regfile_5; // @[registerFile.scala 25:26]
  reg [31:0] reg_regfile_6; // @[registerFile.scala 25:26]
  reg [31:0] reg_regfile_7; // @[registerFile.scala 25:26]
  reg [31:0] reg_regfile_8; // @[registerFile.scala 25:26]
  reg [31:0] reg_regfile_9; // @[registerFile.scala 25:26]
  reg [31:0] reg_regfile_10; // @[registerFile.scala 25:26]
  reg [31:0] reg_regfile_11; // @[registerFile.scala 25:26]
  reg [31:0] reg_regfile_12; // @[registerFile.scala 25:26]
  reg [31:0] reg_regfile_13; // @[registerFile.scala 25:26]
  reg [31:0] reg_regfile_14; // @[registerFile.scala 25:26]
  reg [31:0] reg_regfile_15; // @[registerFile.scala 25:26]
  reg [31:0] reg_regfile_16; // @[registerFile.scala 25:26]
  reg [31:0] reg_regfile_17; // @[registerFile.scala 25:26]
  reg [31:0] reg_regfile_18; // @[registerFile.scala 25:26]
  reg [31:0] reg_regfile_19; // @[registerFile.scala 25:26]
  reg [31:0] reg_regfile_20; // @[registerFile.scala 25:26]
  reg [31:0] reg_regfile_21; // @[registerFile.scala 25:26]
  reg [31:0] reg_regfile_22; // @[registerFile.scala 25:26]
  reg [31:0] reg_regfile_23; // @[registerFile.scala 25:26]
  reg [31:0] reg_regfile_24; // @[registerFile.scala 25:26]
  reg [31:0] reg_regfile_25; // @[registerFile.scala 25:26]
  reg [31:0] reg_regfile_26; // @[registerFile.scala 25:26]
  reg [31:0] reg_regfile_27; // @[registerFile.scala 25:26]
  reg [31:0] reg_regfile_28; // @[registerFile.scala 25:26]
  reg [31:0] reg_regfile_29; // @[registerFile.scala 25:26]
  reg [31:0] reg_regfile_30; // @[registerFile.scala 25:26]
  reg [31:0] reg_regfile_31; // @[registerFile.scala 25:26]
  wire [31:0] _GEN_65 = 5'h1 == io_b_rport_0_addr ? reg_regfile_1 : reg_regfile_0; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_66 = 5'h2 == io_b_rport_0_addr ? reg_regfile_2 : _GEN_65; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_67 = 5'h3 == io_b_rport_0_addr ? reg_regfile_3 : _GEN_66; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_68 = 5'h4 == io_b_rport_0_addr ? reg_regfile_4 : _GEN_67; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_69 = 5'h5 == io_b_rport_0_addr ? reg_regfile_5 : _GEN_68; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_70 = 5'h6 == io_b_rport_0_addr ? reg_regfile_6 : _GEN_69; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_71 = 5'h7 == io_b_rport_0_addr ? reg_regfile_7 : _GEN_70; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_72 = 5'h8 == io_b_rport_0_addr ? reg_regfile_8 : _GEN_71; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_73 = 5'h9 == io_b_rport_0_addr ? reg_regfile_9 : _GEN_72; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_74 = 5'ha == io_b_rport_0_addr ? reg_regfile_10 : _GEN_73; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_75 = 5'hb == io_b_rport_0_addr ? reg_regfile_11 : _GEN_74; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_76 = 5'hc == io_b_rport_0_addr ? reg_regfile_12 : _GEN_75; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_77 = 5'hd == io_b_rport_0_addr ? reg_regfile_13 : _GEN_76; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_78 = 5'he == io_b_rport_0_addr ? reg_regfile_14 : _GEN_77; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_79 = 5'hf == io_b_rport_0_addr ? reg_regfile_15 : _GEN_78; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_80 = 5'h10 == io_b_rport_0_addr ? reg_regfile_16 : _GEN_79; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_81 = 5'h11 == io_b_rport_0_addr ? reg_regfile_17 : _GEN_80; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_82 = 5'h12 == io_b_rport_0_addr ? reg_regfile_18 : _GEN_81; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_83 = 5'h13 == io_b_rport_0_addr ? reg_regfile_19 : _GEN_82; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_84 = 5'h14 == io_b_rport_0_addr ? reg_regfile_20 : _GEN_83; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_85 = 5'h15 == io_b_rport_0_addr ? reg_regfile_21 : _GEN_84; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_86 = 5'h16 == io_b_rport_0_addr ? reg_regfile_22 : _GEN_85; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_87 = 5'h17 == io_b_rport_0_addr ? reg_regfile_23 : _GEN_86; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_88 = 5'h18 == io_b_rport_0_addr ? reg_regfile_24 : _GEN_87; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_89 = 5'h19 == io_b_rport_0_addr ? reg_regfile_25 : _GEN_88; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_90 = 5'h1a == io_b_rport_0_addr ? reg_regfile_26 : _GEN_89; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_91 = 5'h1b == io_b_rport_0_addr ? reg_regfile_27 : _GEN_90; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_92 = 5'h1c == io_b_rport_0_addr ? reg_regfile_28 : _GEN_91; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_93 = 5'h1d == io_b_rport_0_addr ? reg_regfile_29 : _GEN_92; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_94 = 5'h1e == io_b_rport_0_addr ? reg_regfile_30 : _GEN_93; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_97 = 5'h1 == io_b_rport_1_addr ? reg_regfile_1 : reg_regfile_0; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_98 = 5'h2 == io_b_rport_1_addr ? reg_regfile_2 : _GEN_97; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_99 = 5'h3 == io_b_rport_1_addr ? reg_regfile_3 : _GEN_98; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_100 = 5'h4 == io_b_rport_1_addr ? reg_regfile_4 : _GEN_99; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_101 = 5'h5 == io_b_rport_1_addr ? reg_regfile_5 : _GEN_100; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_102 = 5'h6 == io_b_rport_1_addr ? reg_regfile_6 : _GEN_101; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_103 = 5'h7 == io_b_rport_1_addr ? reg_regfile_7 : _GEN_102; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_104 = 5'h8 == io_b_rport_1_addr ? reg_regfile_8 : _GEN_103; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_105 = 5'h9 == io_b_rport_1_addr ? reg_regfile_9 : _GEN_104; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_106 = 5'ha == io_b_rport_1_addr ? reg_regfile_10 : _GEN_105; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_107 = 5'hb == io_b_rport_1_addr ? reg_regfile_11 : _GEN_106; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_108 = 5'hc == io_b_rport_1_addr ? reg_regfile_12 : _GEN_107; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_109 = 5'hd == io_b_rport_1_addr ? reg_regfile_13 : _GEN_108; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_110 = 5'he == io_b_rport_1_addr ? reg_regfile_14 : _GEN_109; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_111 = 5'hf == io_b_rport_1_addr ? reg_regfile_15 : _GEN_110; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_112 = 5'h10 == io_b_rport_1_addr ? reg_regfile_16 : _GEN_111; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_113 = 5'h11 == io_b_rport_1_addr ? reg_regfile_17 : _GEN_112; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_114 = 5'h12 == io_b_rport_1_addr ? reg_regfile_18 : _GEN_113; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_115 = 5'h13 == io_b_rport_1_addr ? reg_regfile_19 : _GEN_114; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_116 = 5'h14 == io_b_rport_1_addr ? reg_regfile_20 : _GEN_115; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_117 = 5'h15 == io_b_rport_1_addr ? reg_regfile_21 : _GEN_116; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_118 = 5'h16 == io_b_rport_1_addr ? reg_regfile_22 : _GEN_117; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_119 = 5'h17 == io_b_rport_1_addr ? reg_regfile_23 : _GEN_118; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_120 = 5'h18 == io_b_rport_1_addr ? reg_regfile_24 : _GEN_119; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_121 = 5'h19 == io_b_rport_1_addr ? reg_regfile_25 : _GEN_120; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_122 = 5'h1a == io_b_rport_1_addr ? reg_regfile_26 : _GEN_121; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_123 = 5'h1b == io_b_rport_1_addr ? reg_regfile_27 : _GEN_122; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_124 = 5'h1c == io_b_rport_1_addr ? reg_regfile_28 : _GEN_123; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_125 = 5'h1d == io_b_rport_1_addr ? reg_regfile_29 : _GEN_124; // @[registerFile.scala 40:28]
  wire [31:0] _GEN_126 = 5'h1e == io_b_rport_1_addr ? reg_regfile_30 : _GEN_125; // @[registerFile.scala 40:28]
  assign io_b_rport_0_data = 5'h1f == io_b_rport_0_addr ? reg_regfile_31 : _GEN_94; // @[registerFile.scala 40:28]
  assign io_b_rport_1_data = 5'h1f == io_b_rport_1_addr ? reg_regfile_31 : _GEN_126; // @[registerFile.scala 40:28]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_regfile_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  reg_regfile_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reg_regfile_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  reg_regfile_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  reg_regfile_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  reg_regfile_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  reg_regfile_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  reg_regfile_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  reg_regfile_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  reg_regfile_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  reg_regfile_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  reg_regfile_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  reg_regfile_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  reg_regfile_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  reg_regfile_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  reg_regfile_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  reg_regfile_16 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  reg_regfile_17 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  reg_regfile_18 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  reg_regfile_19 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  reg_regfile_20 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  reg_regfile_21 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  reg_regfile_22 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  reg_regfile_23 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  reg_regfile_24 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  reg_regfile_25 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  reg_regfile_26 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  reg_regfile_27 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  reg_regfile_28 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  reg_regfile_29 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  reg_regfile_30 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  reg_regfile_31 = _RAND_31[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (io_b_wport_0_en) begin
      if (5'h0 == io_b_wport_0_addr) begin
        reg_regfile_0 <= io_b_wport_0_data;
      end
    end
    if (io_b_wport_0_en) begin
      if (5'h1 == io_b_wport_0_addr) begin
        reg_regfile_1 <= io_b_wport_0_data;
      end
    end
    if (io_b_wport_0_en) begin
      if (5'h2 == io_b_wport_0_addr) begin
        reg_regfile_2 <= io_b_wport_0_data;
      end
    end
    if (io_b_wport_0_en) begin
      if (5'h3 == io_b_wport_0_addr) begin
        reg_regfile_3 <= io_b_wport_0_data;
      end
    end
    if (io_b_wport_0_en) begin
      if (5'h4 == io_b_wport_0_addr) begin
        reg_regfile_4 <= io_b_wport_0_data;
      end
    end
    if (io_b_wport_0_en) begin
      if (5'h5 == io_b_wport_0_addr) begin
        reg_regfile_5 <= io_b_wport_0_data;
      end
    end
    if (io_b_wport_0_en) begin
      if (5'h6 == io_b_wport_0_addr) begin
        reg_regfile_6 <= io_b_wport_0_data;
      end
    end
    if (io_b_wport_0_en) begin
      if (5'h7 == io_b_wport_0_addr) begin
        reg_regfile_7 <= io_b_wport_0_data;
      end
    end
    if (io_b_wport_0_en) begin
      if (5'h8 == io_b_wport_0_addr) begin
        reg_regfile_8 <= io_b_wport_0_data;
      end
    end
    if (io_b_wport_0_en) begin
      if (5'h9 == io_b_wport_0_addr) begin
        reg_regfile_9 <= io_b_wport_0_data;
      end
    end
    if (io_b_wport_0_en) begin
      if (5'ha == io_b_wport_0_addr) begin
        reg_regfile_10 <= io_b_wport_0_data;
      end
    end
    if (io_b_wport_0_en) begin
      if (5'hb == io_b_wport_0_addr) begin
        reg_regfile_11 <= io_b_wport_0_data;
      end
    end
    if (io_b_wport_0_en) begin
      if (5'hc == io_b_wport_0_addr) begin
        reg_regfile_12 <= io_b_wport_0_data;
      end
    end
    if (io_b_wport_0_en) begin
      if (5'hd == io_b_wport_0_addr) begin
        reg_regfile_13 <= io_b_wport_0_data;
      end
    end
    if (io_b_wport_0_en) begin
      if (5'he == io_b_wport_0_addr) begin
        reg_regfile_14 <= io_b_wport_0_data;
      end
    end
    if (io_b_wport_0_en) begin
      if (5'hf == io_b_wport_0_addr) begin
        reg_regfile_15 <= io_b_wport_0_data;
      end
    end
    if (io_b_wport_0_en) begin
      if (5'h10 == io_b_wport_0_addr) begin
        reg_regfile_16 <= io_b_wport_0_data;
      end
    end
    if (io_b_wport_0_en) begin
      if (5'h11 == io_b_wport_0_addr) begin
        reg_regfile_17 <= io_b_wport_0_data;
      end
    end
    if (io_b_wport_0_en) begin
      if (5'h12 == io_b_wport_0_addr) begin
        reg_regfile_18 <= io_b_wport_0_data;
      end
    end
    if (io_b_wport_0_en) begin
      if (5'h13 == io_b_wport_0_addr) begin
        reg_regfile_19 <= io_b_wport_0_data;
      end
    end
    if (io_b_wport_0_en) begin
      if (5'h14 == io_b_wport_0_addr) begin
        reg_regfile_20 <= io_b_wport_0_data;
      end
    end
    if (io_b_wport_0_en) begin
      if (5'h15 == io_b_wport_0_addr) begin
        reg_regfile_21 <= io_b_wport_0_data;
      end
    end
    if (io_b_wport_0_en) begin
      if (5'h16 == io_b_wport_0_addr) begin
        reg_regfile_22 <= io_b_wport_0_data;
      end
    end
    if (io_b_wport_0_en) begin
      if (5'h17 == io_b_wport_0_addr) begin
        reg_regfile_23 <= io_b_wport_0_data;
      end
    end
    if (io_b_wport_0_en) begin
      if (5'h18 == io_b_wport_0_addr) begin
        reg_regfile_24 <= io_b_wport_0_data;
      end
    end
    if (io_b_wport_0_en) begin
      if (5'h19 == io_b_wport_0_addr) begin
        reg_regfile_25 <= io_b_wport_0_data;
      end
    end
    if (io_b_wport_0_en) begin
      if (5'h1a == io_b_wport_0_addr) begin
        reg_regfile_26 <= io_b_wport_0_data;
      end
    end
    if (io_b_wport_0_en) begin
      if (5'h1b == io_b_wport_0_addr) begin
        reg_regfile_27 <= io_b_wport_0_data;
      end
    end
    if (io_b_wport_0_en) begin
      if (5'h1c == io_b_wport_0_addr) begin
        reg_regfile_28 <= io_b_wport_0_data;
      end
    end
    if (io_b_wport_0_en) begin
      if (5'h1d == io_b_wport_0_addr) begin
        reg_regfile_29 <= io_b_wport_0_data;
      end
    end
    if (io_b_wport_0_en) begin
      if (5'h1e == io_b_wport_0_addr) begin
        reg_regfile_30 <= io_b_wport_0_data;
      end
    end
    if (io_b_wport_0_en) begin
      if (5'h1f == io_b_wport_0_addr) begin
        reg_regfile_31 <= io_b_wport_0_data;
      end
    end
  end
endmodule
